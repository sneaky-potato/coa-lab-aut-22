`timescale 1ns / 1ps

/*
/////////////////////////////////////////////
//// COA LAB Assignment 6                ////
//// Group Number 23                     ////
//// Ashwani Kumar Kamal (20CS10011)     ////
//// Astitva (20CS30007)                 ////
/////////////////////////////////////////////
*/

// ALU module to compute the result and flags based on ALUop and ALUsel

module ALU (
    input signed [31:0] in1, 
    input signed [31:0] in2, 
    input ALUsel, 
    input [4:0] ALUop, 
    output reg carry,
    output reg zero, 
    output reg sign, 
    output reg [31:0] result
    );

    // Stores carry generated by adder1
    wire carryTemp;

    // Stores 32-bit output of not, adder1, shifter, and, xor, mux1, mux2 respectively from left to right.
    wire [31:0] not1Out, adder1Out, shifterOut, and1Out, xor1Out, mux1Out, mux2Out;

    mux_32b_2_1 mux1 (.in1(a), .in2(32'd1), .sel(ALUsel), .out(mux1Out));
    mux_32b_2_1 mux2 (.in1(b), .in2(not1Out), .sel(ALUsel), .out(mux2Out));

    cla_32_lcu adder1(.in1(mux1Out), .in2(mux2Out), .cin(1'b0), .cout(carryTemp), .out(adder1Out));

    shifter shifter1 (.in(mux1Out), .shamt(mux2Out), .left_shift(ALUop[1]), .out(shifterOut), .arithmetic_shift(ALUop[0]));

    assign not1Out = ~b;
    assign and1Out = mux1Out & mux2Out;
    assign xor1Out = mux1Out ^ mux2Out;

    // result changes on change of any input signal
    always @(*) begin
        if (ALUop == 5'b00000) begin
            result = mux1Out;
        end else if (ALUop == 5'b00001) begin
            carry = carryTemp;
            result = adder1Out;
        end else if (ALUop == 5'b00101) begin
            result = adder1Out;
        end else if (ALUop == 5'b10101) begin
            result = adder1Out;
        end else if (ALUop == 5'b00010) begin
            result = and1Out;
        end else if (ALUop == 5'b00011) begin
            result = xor1Out;
        end else if (ALUop[4:2] == 3'b010) begin
            result = shifterOut;
        end 
        else begin
            result = 32'd0;
        end
    end

    // Flags change on change of result
    always @(result) begin
        if (!result) begin
            zero = 1'b1;
        end else begin
            zero = 1'b0;
        end
        sign = result[31];
    end
    
endmodule
